`timescale 1ns/10ps
`include "adder_64.v"

module adder_test;

reg signed [63:0] a;
reg signed [63:0] b;


wire signed [63:0] sum;
wire overflow, carry;

adder_64 tt(
.a(a),
.b(b),
.sum(sum),
.overflow(overflow),
.carry(carry));




initial begin

    $dumpfile("test.vcd");
    $dumpvars(0,adder_test);
   
     a = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    b = 64'b1111111111111111111111111111111111111111111111111111111111111111;

    #5;
    
    a = 64'b1111111111111111111111111111111111111111111111111111111111111101;
    b = 64'b1111111111111111111111111111111111111111111111111111111111110111;

    #5;

    a = 64'b1111111111111111111111111111111111101111111111111111111111111110;
    b = 64'b1111111111111111111111111111111111011111111111111111111111111101;

    #5;

    
    a = 64'b0111111111111111111111111111111111111111111111111111111111111111;
    b = 64'b0111111111111111111111111111111111111111111111111111111111111111;
    #5;

    a = 64'b1000000000000000000000000000000000000000000000000000000000000001;
    b = 64'b1000000000000000000000000000000000000000000000000000000000000001;
    #5;
end
  
endmodule

