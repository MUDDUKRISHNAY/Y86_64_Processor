`timescale 1ns/10ps
`include "subtractor_64.v"

module subtractor_test;

    reg signed [63:0] a;
    reg signed [63:0] b;
    

    wire signed [63:0] difference;
    wire overflow, borrow;

    subtractor_64 sub (
        .a(a),
        .b(b),
        .difference(difference),
        .overflow(overflow),
        .borrow(borrow)
    );

    
    initial begin
        $dumpfile("test.vcd");
        $dumpvars(0, subtractor_test);
        

        a = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        b = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        #8;

        a = 64'b1111111111111111111111111111111111111111111111111111111111111110;
        b = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        #8;

        a = 64'b1111111111111111111111111111111111111111111111111111111111111101;
        b = 64'b1111111111111111111111111111111111111111111111111111111111111110;
        #8;

        a = 64'b1111111111111111111111111111111111111111111111111111111111111100;
        b = 64'b1111111111111111111111111111111111111111111111111111111111111101;
        #10;

        a = 64'b1111111111111111111111111111111111111111111111111111111111111011;
        b = 64'b1111111111111111111111111111111111111111111111111111111111111100;
        #10;

        a = 64'b0111111111111111111111111111111111111111111111111111111111111111;
        b = 64'b1111111111111111111111111111111111111111111111111111111111100001;
        #10;

        a = 64'b0110010111100000000000000111111111110000110101010101010100000000;
        b = 64'b0111111100000000000000000000000000000000000000000000000001010101;
        #10;
    end


endmodule

