`timescale 1ns/10ps
`include "AND.v"

module and_tb;

    reg signed [63:0] a;
    reg signed [63:0] b;
    wire signed [63:0] ans;

    and_64 andi(a, b, ans);

    initial begin
        $dumpfile("test.vcd");
        $dumpvars(0, and_tb);

        a= 64'b1111111111111111111111111111111111111111111111111111111111111111;
        b = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        #10;

        a = 64'b1111111111111111111111111111111111111111111111111111111111111110;
        b = 64'b1111111111111111111111111111111111111111111111111111111111111110;
        #10;

        a = 64'b1111111111111111111111111111111111111111111111111111111111111101;
        b = 64'b1111111111111111111111111111111111111111111111111111111111111101;
        #10;

        a = 64'b1111111111111111111111111111111111111111111111111111111111111100;
        b = 64'b1111111111111111111111111111111111111111111111111111111111111100;
        #10;

        a = 64'b1111111111111111111111111111111111111111111111111111111111111011;
        b = 64'b1111111111111111111111111111111111111111111111111111111111111011;
        #10;

        a = 64'b0000000000000000000000000000000000000000000000000000000000000001;
        b = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        #10;

        a = 64'b1010101010101010101010101010101010101010101010101010101010101010;
        b = 64'b0101010101010101010101010101010101010101010101010101010101010101;
        #10;

        a = 64'b1111000011110000111100001111000011110000111100001111000011110000;
        b = 64'b0000111100001111000011110000111100001111000011110000111100001111;
        #10;

        a = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        b = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        #10;

        a = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        b = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        #10;
    end

endmodule
